----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:02:17 11/11/2014 
-- Design Name: 
-- Module Name:    ffD_reset - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ffD_reset is
    Port ( d : in  STD_LOGIC_VECTOR(3 downto 0);
           clk : in  STD_LOGIC;
           ce : in  STD_LOGIC;
           q : out  STD_LOGIC_VECTOR(3 downto 0);
           reset : in  STD_LOGIC
			  );
end ffD_reset;

architecture Behavioral of ffD_reset is

begin

process(clk,reset)

begin

	if reset='1' then
			q<= "0000";
	elsif (clk'event and clk='1') then
		if ce= '1' then
			q <= d;
			end if;
		end if;
			
end process;
		



end Behavioral;

